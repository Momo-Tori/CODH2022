module decoder_4t16 (
    input[3:0] i,
    output reg[15:0] o
);
always @(*) begin
    case (i)
        0:o=16'b1;
        1:o=16'b10;
        2:o=16'b100;
        3:o=16'b1000;
        4:o=16'b10000;
        5:o=16'b100000;
        6:o=16'b1000000;
        7:o=16'b10000000;
        8:o=16'b100000000;
        9:o=16'b1000000000;
       10:o=16'b10000000000;
       11:o=16'b100000000000;
       12:o=16'b1000000000000;
       13:o=16'b10000000000000;
       14:o=16'b100000000000000;
       15:o=16'b1000000000000000;
    endcase
end
endmodule //decoder