`timescale 1ns / 1ps
module tb( );
reg [5:0] a;
reg [5:0]b;
reg [2:0]s;
wire [5:0] y;     //运算结果
wire [2:0] f;
initial
begin
a=0;b=0;
begin
#5 a=6'b100000;b=6'b100000;//s=0
#5 a=6'b101100;b=6'b011111;
#5 a=6'b001100;b=6'b100000;
#5 a=6'b001010;b=6'b001010;
#5 a=6'b011001;b=6'b011111;
#5 a=6'b011111;b=6'b000001;
#5 a=6'b011111; b=6'b100000;
#5 a=6'b000001; b=6'b111111;

#5 a=6'b100000;b=6'b100000;//s=1
#5 a=6'b101100;b=6'b011111;
#5 a=6'b001100;b=6'b100000;
#5 a=6'b001010;b=6'b001010;
#5 a=6'b011001;b=6'b011111;
#5 a=6'b011111;b=6'b000001;
#5 a=6'b011111; b=6'b100000;
#5 a=6'b000001; b=6'b111111;

#5 a=6'b100000;b=6'b100000;//s=2
#5 a=6'b101100;b=6'b011111;
#5 a=6'b001100;b=6'b100000;
#5 a=6'b001010;b=6'b001010;
#5 a=6'b011001;b=6'b011111;
#5 a=6'b011111;b=6'b000001;
#5 a=6'b011111; b=6'b100000;
#5 a=6'b000001; b=6'b111111;

#5 a=6'b100000;b=6'b100000;//s=3
#5 a=6'b101100;b=6'b011111;
#5 a=6'b001100;b=6'b100000;
#5 a=6'b001010;b=6'b001010;
#5 a=6'b011001;b=6'b011111;
#5 a=6'b011111;b=6'b000001;
#5 a=6'b011111; b=6'b100000;
#5 a=6'b000001; b=6'b111111;

#5 a=6'b100000;b=6'b100000;//s=4
#5 a=6'b101100;b=6'b011111;
#5 a=6'b001100;b=6'b100000;
#5 a=6'b001010;b=6'b001010;
#5 a=6'b011001;b=6'b011111;
#5 a=6'b011111;b=6'b000001;
#5 a=6'b011111; b=6'b100000;
#5 a=6'b000001; b=6'b111111;

#5 a=6'b100000;b=6'b000011;//s=5
#5 a=6'b101100;b=6'b000011;
#5 a=6'b001100;b=6'b000010;
#5 a=6'b001010;b=6'b000001;
#5 a=6'b011001;b=6'b011111;
#5 a=6'b011111;b=6'b000001;
#5 a=6'b011111; b=6'b000010;
#5 a=6'b000001; b=6'b000001;

#5 a=6'b100000;b=6'b000011;//s=6
#5 a=6'b101100;b=6'b000011;
#5 a=6'b001100;b=6'b000010;
#5 a=6'b001010;b=6'b000001;
#5 a=6'b011001;b=6'b011111;
#5 a=6'b011111;b=6'b000001;
#5 a=6'b011111; b=6'b000010;
#5 a=6'b000001; b=6'b000001;

#5 a=6'b100000;b=6'b000011;//s=7
#5 a=6'b101100;b=6'b000011;
#5 a=6'b001100;b=6'b000010;
#5 a=6'b001010;b=6'b000001;
#5 a=6'b011001;b=6'b011111;
#5 a=6'b011111;b=6'b000001;
#5 a=6'b011111; b=6'b000010;
#5 a=6'b000001; b=6'b000001;
end
end

initial
begin
s=0;
forever
#40 s=s+1;
end
initial
#320 $stop;

alu#(6) alu(
.a(a),
.b(b),
.s(s),
.y(y),
.f(f));
endmodule